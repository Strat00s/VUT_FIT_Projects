-- fsm.vhd: Finite State Machine
-- Author(s): 
--
library ieee;
use ieee.std_logic_1164.all;
-- ----------------------------------------------------------------------------
--                        Entity declaration
-- ----------------------------------------------------------------------------
entity fsm is
port(
   CLK         : in  std_logic;
   RESET       : in  std_logic;

   -- Input signals
   KEY         : in  std_logic_vector(15 downto 0);
   CNT_OF      : in  std_logic;

   -- Output signals
   FSM_CNT_CE  : out std_logic;
   FSM_MX_MEM  : out std_logic;
   FSM_MX_LCD  : out std_logic;
   FSM_LCD_WR  : out std_logic;
   FSM_LCD_CLR : out std_logic
);
end entity fsm;

-- ----------------------------------------------------------------------------
--                      Architecture declaration
-- ----------------------------------------------------------------------------
architecture behavioral of fsm is
	-- xbasty00 : kod1 = 1063475812 	 kod2 = 1065026509
   type t_state is (K_1, K_10, K_106, K_1063, K_10634, K_106347, K_1063475, K_10634758, K_106347581, K_1063475812,
												  K_1065, K_10650, K_106502, K_1065026, K_10650265, K_106502650, K_1065026509,
						  DEFAULT, ERROR, MSG_ERROR, MSG_OK, FINISH);
   signal present_state, next_state : t_state;

begin
-- -------------------------------------------------------
sync_logic : process(RESET, CLK)
begin
   if (RESET = '1') then
      present_state <= DEFAULT;
   elsif (CLK'event AND CLK = '1') then
      present_state <= next_state;
   end if;
end process sync_logic;

-- -------------------------------------------------------
-- -------------------------------------------------------
-- -------------------------------------------------------
next_state_logic : process(present_state, KEY, CNT_OF)
begin
   case (present_state) is
	-- key preses
   -- - - - - - - - - - - - - - - - - - - - - - -
	-- start
   when DEFAULT =>
      next_state <= DEFAULT;
		if (KEY(1) = '1') then
			next_state <= K_1;
      elsif (KEY(15) = '1') then			-- when # is pressed, got to error
         next_state <= MSG_ERROR;
      elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= ERROR;
      end if;
	
	-- wrong key
	-- once any wrong key was pressed, just loop here till # is pressed and then print error msg
	when ERROR =>
      next_state <= ERROR;
      if (KEY(15) = '1') then			-- when # is pressed, got to error
         next_state <= MSG_ERROR;
      end if;
	
	--	1
   when K_1 =>
      next_state <= K_1;
		if (KEY(0) = '1') then
			next_state <= K_10;
      elsif (KEY(15) = '1') then			-- when # is pressed, got to error
         next_state <= MSG_ERROR;
      elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= ERROR;
      end if;
		
	-- 10	
	when K_10 =>
      next_state <= K_10;
		if (KEY(6) = '1') then
			next_state <= K_106;
      elsif (KEY(15) = '1') then			-- when # is pressed, got to error
         next_state <= MSG_ERROR;
      elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= ERROR;
      end if;
	
	-- 106
	when K_106 =>
      next_state <= K_106;
		if (KEY(3) = '1') then
			next_state <= K_1063;
		elsif (KEY(5) = '1') then		-- TODO check if this works 
			next_state <= K_1065;
      elsif (KEY(15) = '1') then
         next_state <= MSG_ERROR;
      elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= ERROR;
      end if;
		
	-- 1063
	when K_1063 =>
      next_state <= K_1063;
		if (KEY(4) = '1') then
			next_state <= K_10634;
      elsif (KEY(15) = '1') then
         next_state <= MSG_ERROR;
      elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= ERROR;
      end if;

	-- 10634
	when K_10634 =>
      next_state <= K_10634;
		if (KEY(7) = '1') then
			next_state <= K_106347;
      elsif (KEY(15) = '1') then
         next_state <= MSG_ERROR;
      elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= ERROR;
      end if;

	-- 106347
	when K_106347 =>
      next_state <= K_106347;
		if (KEY(5) = '1') then
			next_state <= K_1063475;
      elsif (KEY(15) = '1') then
         next_state <= MSG_ERROR;
      elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= ERROR;
      end if;
		
	-- 1063475
	when K_1063475 =>
      next_state <= K_1063475;
		if (KEY(8) = '1') then
			next_state <= K_10634758;
      elsif (KEY(15) = '1') then
         next_state <= MSG_ERROR;
      elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= ERROR;
      end if;
		
	-- 10634758
	when K_10634758 =>
      next_state <= K_10634758;
		if (KEY(1) = '1') then
			next_state <= K_106347581;
      elsif (KEY(15) = '1') then
         next_state <= MSG_ERROR;
      elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= ERROR;
      end if;
		
	-- 106347581
	when K_106347581 =>
      next_state <= K_106347581;
		if (KEY(2) = '1') then
			next_state <= K_1063475812;
      elsif (KEY(15) = '1') then
         next_state <= MSG_ERROR;
      elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= ERROR;
      end if;
		
	-- 1063475812
	when K_1063475812 =>
      next_state <= K_1063475812;
      if (KEY(15) = '1') then
         next_state <= MSG_OK;		-- end of code, go print OK message
      elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= ERROR;
      end if;
		
	-- 1065	
	when K_1065 =>
      next_state <= K_1065;
		if (KEY(0) = '1') then
			next_state <= K_10650;
      elsif (KEY(15) = '1') then			-- when # is pressed, got to error
         next_state <= MSG_ERROR;
      elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= ERROR;
      end if;

	-- 10650
	when K_10650 =>
      next_state <= K_10650;
		if (KEY(2) = '1') then
			next_state <= K_106502;
      elsif (KEY(15) = '1') then			-- when # is pressed, got to error
         next_state <= MSG_ERROR;
      elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= ERROR;
      end if;
		
	-- 106502
	when K_106502 =>
      next_state <= K_106502;
		if (KEY(6) = '1') then
			next_state <= K_1065026;
      elsif (KEY(15) = '1') then			-- when # is pressed, got to error
         next_state <= MSG_ERROR;
      elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= ERROR;
      end if;
		
	-- 1065026
	when K_1065026 =>
      next_state <= K_1065026;
		if (KEY(5) = '1') then
			next_state <= K_10650265;
      elsif (KEY(15) = '1') then			-- when # is pressed, got to error
         next_state <= MSG_ERROR;
      elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= ERROR;
      end if;
		
	-- 10650265
	when K_10650265 =>
      next_state <= K_10650265;
		if (KEY(0) = '1') then
			next_state <= K_106502650;
      elsif (KEY(15) = '1') then			-- when # is pressed, got to error
         next_state <= MSG_ERROR;
      elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= ERROR;
      end if;

	-- 106502650
	when K_106502650 =>
      next_state <= K_106502650;
		if (KEY(9) = '1') then
			next_state <= K_1065026509;
      elsif (KEY(15) = '1') then			-- when # is pressed, got to error
         next_state <= MSG_ERROR;
      elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= ERROR;
      end if;

	-- 1065026509
	when K_1065026509 =>
      next_state <= K_1065026509;
		if (KEY(15) = '1') then
         next_state <= MSG_OK;		-- end of code, go print OK message
      elsif (KEY(14 downto 0) /= "000000000000000") then
			next_state <= ERROR;
      end if;

	-- MESSAGES
   -- - - - - - - - - - - - - - - - - - - - - - -
   when MSG_ERROR =>
      next_state <= MSG_ERROR;
      if (CNT_OF = '1') then
         next_state <= FINISH;
      end if;
   -- - - - - - - - - - - - - - - - - - - - - - -
   when MSG_OK =>
      next_state <= MSG_OK;
      if (CNT_OF = '1') then
         next_state <= FINISH;
      end if;
   -- - - - - - - - - - - - - - - - - - - - - - -
	
   when FINISH =>
      next_state <= FINISH;
      if (KEY(15) = '1') then
         next_state <= DEFAULT; 
      end if;
   -- - - - - - - - - - - - - - - - - - - - - - -
   when others =>
      next_state <= DEFAULT;
   end case;
end process next_state_logic;

-- -------------------------------------------------------
output_logic : process(present_state, KEY)
begin
   FSM_CNT_CE     <= '0';
   FSM_MX_MEM     <= '0';
   FSM_MX_LCD     <= '0';
   FSM_LCD_WR     <= '0';
   FSM_LCD_CLR    <= '0';

   case (present_state) is
   -- - - - - - - - - - - - - - - - - - - - - - -
	-- print *
   when DEFAULT | ERROR | K_1 | K_10 | K_106 | K_1063 | K_10634 | K_106347 | K_1063475 | K_10634758 | K_106347581 | K_1063475812 |
													K_1065 | K_10650 | K_106502 | K_1065026 | K_10650265 | K_106502650 | K_1065026509 =>	-- add allt states to print *
      if (KEY(14 downto 0) /= "000000000000000") then
         FSM_LCD_WR     <= '1';
      end if;
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
   -- - - - - - - - - - - - - - - - - - - - - - -
   when MSG_ERROR =>
      FSM_CNT_CE     <= '1';
      FSM_MX_LCD     <= '1';
      FSM_LCD_WR     <= '1';
   -- - - - - - - - - - - - - - - - - - - - - - -
   when MSG_OK =>
      FSM_CNT_CE     <= '1';
      FSM_MX_LCD     <= '1';
      FSM_LCD_WR     <= '1';
		FSM_MX_MEM		<= '1';	-- print pritstup povolen
   -- - - - - - - - - - - - - - - - - - - - - - -
   when FINISH =>
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
   -- - - - - - - - - - - - - - - - - - - - - - -
   when others =>
   end case;
end process output_logic;

end architecture behavioral;

